/*
 * WIP floating point unit
 * Should end up supporting FP16, FP32, and FP64
 */
