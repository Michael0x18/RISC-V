`default_nettype none
module decode(
	input wire[31:0] instruction
//TODO others
);


endmodule /*decode*/
`default_nettype wire
